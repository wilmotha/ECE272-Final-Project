module math(input logic [5:0] num1
			input)