module LED_top_module( 
	/**************************/
	/* Set inputs and outputs */
	/* to the whole FPGA here */
	/**************************/
	input logic [7:0] button,
	input logic reset_n,
	output logic [6:0] sevenseg,
	output logic [2:0] state
	);
		/*******************************/
		/* Set internal variables here */
		/*******************************/
		logic clk;		//used for the oscillator's 2.08 MHz clock
		logic clk_slow;	//used for slowed down, 5 Hz clock
		logic clk_manual = 1'b1; //Initialize the manual clock to start
		logic clk_manual_memory;
		
		logic [2:0] num_state; 	//look at Operation_State_Machine to understand this
		logic [2:0] adr;			//Adress in the memory
		
		logic [3:0] thous;
		logic [3:0] hundr;
		logic [3:0] tens;
		logic [3:0] ones;
		
		logic [3:0] muxToDec;
		
		/***********************/
		/* Define modules here */
		/***********************/
		/*
		parser in( .b(button),
					.thous(thous),
					.hunds(hundr),
					.tens(tens),
					.ones(ones));
		
		mux4 which( .thous(thous),
						.hundr(hundr),
						.tens(tens),
						.ones(ones),
						.s(state),
						.y(muxToDec));
						
		decoder fin( .data(muxToDec),
							.segments(sevenseg)); */
		
		//This is an instance of a special, built in module that accesses our chip's oscillator
		OSCH #("2.08") osc_int (	//"2.08" specifies the operating frequency, 2.08 MHz.
									//Other clock frequencies can be found in the MachX02's documentation
			.STDBY(1'b0),			//Specifies active state
			.OSC(clk),				//Outputs clock signal to 'clk' net
			.SEDSTDBY());			//Leaves SEDSTDBY pin unconnected
		
		
		//This module is instantiated from another file, 'Clock_Counter.sv'
		//It will take an input clock, slow it down based on parameters set inside of the module, and
		//output the new clock. Reset functionality is also built-in
		clock_counter counter_1(
			.clk_i(clk),
			.reset_n(reset_n),
			.clk_o(clk_slow));
			
		//This module is instantiated from another file, 'State_Machine.sv'
		//It contains a Moore state machine that will take a clock and reset, and output a state
		state_machine FSM_1(
			.clk_i(clk_slow),
			.reset_n(reset_n),
			.state(state));
			
		/************************************************/
		/* Add modules for:								*/
		/* Parser 		Determines the 1000's, 100's,   */
		/*				10's and 1's place of the number*/
		/* Multiplexer	Determines which parser output  */
		/*				to pass to the decoder			*/
		/* Decoder		Convert 4-bit binary to 7-seg   */
		/*				output for numbers 0-9			*/
		/************************************************/
endmodule
